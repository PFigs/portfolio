-----------------------------------------------------------------------------
-- Vhdl model created by vec2mem, (c) 2006-2011 Horacio Neto, Paulo Flores.
-- Command: vec2mem rnd   1073741823 1301579652 
-----------------------------------------------------------------------------

library ieee;
library UNISIM;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use UNISIM.Vcomponents.all;

entity memsdata is
  port ( 
         addrA : in  std_logic_vector(8 downto 0);
         addrB : in  std_logic_vector(8 downto 0);
         addrC : in  std_logic_vector(8 downto 0);
         addrD : in  std_logic_vector(8 downto 0);
         addrE : in  std_logic_vector(8 downto 0);
         addrF : in  std_logic_vector(8 downto 0);
         doA   : out std_logic_vector(31 downto 0);
         doB   : out std_logic_vector(31 downto 0);
         doC   : out std_logic_vector(31 downto 0);
         doD   : out std_logic_vector(31 downto 0);
         doE   : out std_logic_vector(31 downto 0);
         doF   : out std_logic_vector(31 downto 0);
         clk  : in  std_logic
       );

end memsdata;

architecture GENERATED of memsdata is


begin


  MEM_A : RAMB16_S36
    generic map (
      INIT_00       =>
      X"049EB7300A964B1D29AC224830E1EBC5D71CBBEC10D103AA1ACC8E862142CFEE",
      INIT_01       =>
      X"35FAA2C8F2760BCD0C2490981AEF41F7F7F117E936565CBADC2D3CB73703F753",
      INIT_02       =>
      X"D21A1A6EFC3939DE30970DB2E110D23F38120437F2A8D2C3F5E201EC1C03BE3B",
      INIT_03       =>
      X"1DC02FB1F42FC025F56551503C7D5FC3D309BF8CEC58A8501217E5EE2E931CB6",
      INIT_04       =>
      X"25B0DD6A05B282CAFF7336BA2EACE617C113CB9A34DCEB9DC500C3CFD031DFD5",
      INIT_05       =>
      X"24312E56EC8A582E1018011FC82D701BF68FB567DDA1F553FC08DF831BA07370",
      INIT_06       =>
      X"FE5D5559F924EFB7D87C6C6A0FCA38A3E70AD54A1C43328D1F332AF1C5FA030B",
      INIT_07       =>
      X"EB14C92C04D1E1CCC596D509DAE2E9572711B21B116714E4257D98072A945258",
      INIT_08       =>
      X"14C277931EF55C5931DB178F3922042339447EEFEC2894C6F9AECD69CA9798D8",
      INIT_09       =>
      X"12A955D5DA429582F7DC85270CAF52CBF611672DCB522CF93C9751ACEDE3F712",
      INIT_0A       =>
      X"399686D1E5373E13F2D91AD6CF02347926D9E8BA39B42B1F3685C80FD70FB018",
      INIT_0B       =>
      X"C6CCC0D81E4E655FE57A1AB83C352800F3399C3320A838EC369E52F7D856B2DD",
      INIT_0C       =>
      X"EA3608C5ED0D63D61F069C203C5211B3184AEC43C0113FC7CA76FA241F28E821",
      INIT_0D       =>
      X"C74BC60D3AF6966B3A8A0574303C15F6E84D409620476FF2F85F90CF1B9DEDCB",
      INIT_0E       =>
      X"FFDA8F3B39A888CBD35CECDAE783DC5FC01201FB2E25AEC734AAC189310FCD82",
      INIT_0F       =>
      X"1EF3C48FCCFD28A7116290CD3FCADC6EC63067D033142B6E1A50C1B7C9FB3FD0" )
    port map (ADDR  => addrA,
              CLK   => clk,
              DI    => x"00000000",
              DIP   => x"0",
              EN    => '1',
              SSR   => '0',
              WE    => '0',
              DO    => doA,
              DOP   => open);

  MEM_B : RAMB16_S36
    generic map (
      INIT_00       =>
      X"07B2F258C261A569244C14A72C15048D182B9CA4F73EB0D2CD0E686E1BD98AF1",
      INIT_01       =>
      X"0E42E850D43381782AF6C9581D331ACECCE7BB6B300032EE22A9155ADCABA576",
      INIT_02       =>
      X"DFB15CE906FFF67B07FD7315D5B61D19C72567400E54EA4AC259303F1FA18AE1",
      INIT_03       =>
      X"27503DA6C10CD5C8F2DEED5FCB76B2B5E219113AE5E1C4B8FA1421E9E24E34CC",
      INIT_04       =>
      X"F94340B633B54CB201DD7FB2DC979B41EC025A5AFF7BDA49F84B869AFFED55CD",
      INIT_05       =>
      X"EE4DD3D80FFC98291A5E7D990EAC48F7C1B9AFD9062AFC2123B57F9FE486950C",
      INIT_06       =>
      X"C89D2A53D21F27D93C733192264EF588326DCAF1F5733B18DE5182731CB7ADD8",
      INIT_07       =>
      X"EACD2FBDE94E43D5EBC311552ADFD9F001FE0630EAB63B8DF800EC91F687537B",
      INIT_08       =>
      X"0F2E32DBF9E973E50A84D6C8EAA79DD0C0A6332F16CF8A1628CA1E1E240E97EE",
      INIT_09       =>
      X"F72A9B77EB347336E0E47ADD1A72ED9F3CE69F5E10E7E2B4C0147006EE3A5667",
      INIT_0A       =>
      X"D3A2335AEE221D2AFBB78E401D1ADFDFE584F2D7E998666720A7AE4DFF35FD4F",
      INIT_0B       =>
      X"28AA01F9C965847E3EEE7D5EC49B6A0B1E9854C115A0398918D858B633B87AD1",
      INIT_0C       =>
      X"18F43BC2218E6C27E339A90CEAB9E55BD260394C2950352720350E9427B89B7C",
      INIT_0D       =>
      X"D290C706F4EBA226C10F4E55135AC9B73DC106B015DADB1FF2764EDBE34E1911",
      INIT_0E       =>
      X"CDF4119E12740FDA2637D706DA3B96CDFED1DC81F815B9DD1E84088D21B6FCA2",
      INIT_0F       =>
      X"CEBB623DEC559BBF35F1EADDE702C6C103AB99C72C8C665FE8144963FF102FBC" )
    port map (ADDR  => addrB,
              CLK   => clk,
              DI    => x"00000000",
              DIP   => x"0",
              EN    => '1',
              SSR   => '0',
              WE    => '0',
              DO    => doB,
              DOP   => open);

  MEM_C : RAMB16_S36
    generic map (
      INIT_00       =>
      X"1C2D930319D51A8DC2AA07AFF8DF79F2C0E0DECBE11B9B89D5A5D0E61626F970",
      INIT_01       =>
      X"D27640A2DB0BE747CEDA3BD8F0BF4400C87B204119EE99B2EFAFF5ACF520568A",
      INIT_02       =>
      X"3869A7E5D58DECD0E3BC2CFCF9597829C799DB3211481D221321A1232D5E4465",
      INIT_03       =>
      X"0E33377CC18E9F5D286ADD6B380C3E0C32D33D20FC1541ACC21A532F0BD0765F",
      INIT_04       =>
      X"1A74991ED31DBB45E8E930D3E5544295F6F028420F141647E2AA3AE63E10AE51",
      INIT_05       =>
      X"2944D534DBCEAB203DFBA0A53BE690CFC9586A7F22EFB95F2D0C54F71899267F",
      INIT_06       =>
      X"1CA36B9DC2E061D6C66C9D36D0D2F53ECA76B9F130DEB0662D16C842111D41C8",
      INIT_07       =>
      X"E5712F3D0EC665EC1105481AE76080ECC0932E700F76A8BDFEF5A382C886F065",
      INIT_08       =>
      X"DF5CD38433785EB22F7F12C306C3AD05D903C5941C61577FDDDA7C3233AF8300",
      INIT_09       =>
      X"E580FA7E01B6CDBC0483E9221463B8B61871F888E8B53E02166818111C8B67BA",
      INIT_0A       =>
      X"01890BBBDF11123FF2D81645F9021B57026DA6A2EFF7B46FF2957E21F19AB164",
      INIT_0B       =>
      X"F33C8616FE9F69EFD0E2A017FF8D0316D92E3AB2021C3A2B2E87BAFC31CDB9C6",
      INIT_0C       =>
      X"270B3BEAD4DD9CD1FFB8AA5CCA7FD4303580C94E0C404BAADB00C16DEEBD1C49",
      INIT_0D       =>
      X"F3B17559D005759FC134022DC216C3F52A847B22FF7D3472FD92DAD3D620C26C",
      INIT_0E       =>
      X"24A2FA18EE54A760D5302E3A32D540522CCB9BA5361F1BFBFFFD2A0EF3C9804E",
      INIT_0F       =>
      X"F0109DEA36817262FC709EB9C15381A10344EC4C3DD134CA3070E18BC3B7E936" )
    port map (ADDR  => addrC,
              CLK   => clk,
              DI    => x"00000000",
              DIP   => x"0",
              EN    => '1',
              SSR   => '0',
              WE    => '0',
              DO    => doC,
              DOP   => open);

  MEM_D : RAMB16_S36
    generic map (
      INIT_00       =>
      X"D89B2AD308FC703FFA6F0408C27A686721F13456E591673702C1BE0B17716026",
      INIT_01       =>
      X"FD77272CEDCA1829D3251B93C9ADA6DE3A18A2D0C31FA5F4C879A4B13801DEDB",
      INIT_02       =>
      X"FCD14B94EA9A800B18976A30F919625E05F785F3EA42C2D0E3E93424132245A1",
      INIT_03       =>
      X"FC4DB3B33A6C6B453697AA4224DC538D0A5BCD5BC01637E0E86BB4D509084BBA",
      INIT_04       =>
      X"126EB55F146EFB86273B58471A6CD684FBD3D0B3DE3EE808DFFDD27CF959684D",
      INIT_05       =>
      X"FDD602ADF6D9CB013A5170582AB3BD0D3962A3D50C87582F178EA17A2FB4FCF8",
      INIT_06       =>
      X"C2BC43BAD425526EEE6808AAF9B3F800175406DAC3CD88A0211C8DD1DE3AA47C",
      INIT_07       =>
      X"042C9CDC37FDC4BE07847C5ACAD3348FFBB0110C0D181115D43B8A4E16D3BD7F",
      INIT_08       =>
      X"2D2D0205D45DDAB7146F69143D78050D01EF2559C0006D8FD63CACC627824ED5",
      INIT_09       =>
      X"397147B91487CA47DD6970DA1B36A33DD6B1C79A268FA5DA20E532E6EBFE0A8E",
      INIT_0A       =>
      X"1D91190FFAF63A6524EAA100C6BD5B91F839F6AB10C54E92185552E73E85FEAB",
      INIT_0B       =>
      X"F71516A80825FCB8D13EEED90F92C7D3C3F95FDCD9412A1BC80E4B7A39262B4D",
      INIT_0C       =>
      X"0893DDE8D220A2B0CD6216B8DC95D35AE4F3A0AC39043C0108266A46E77B9B9F",
      INIT_0D       =>
      X"D49FB80E02EF3493F3CD6FC9D619B964097DECDA1F45A58238B0488A2E47499D",
      INIT_0E       =>
      X"31C54F713071374FC7CFE91D389F2424D2E01E400CD9AEB9D3B48325CC22C2AF",
      INIT_0F       =>
      X"026CEBE0D6861312FDE4AC05DAF150421F70FC6A35BEAF4DC9B26169CFDE3497" )
    port map (ADDR  => addrD,
              CLK   => clk,
              DI    => x"00000000",
              DIP   => x"0",
              EN    => '1',
              SSR   => '0',
              WE    => '0',
              DO    => doD,
              DOP   => open);

  MEM_E : RAMB16_S36
    generic map (
      INIT_00       =>
      X"CB33AF672B34C78C39812F3CDCEC65CAE2A0E9A527608C8CCF8A4F12C60B164B",
      INIT_01       =>
      X"CA6A9F85DCEAE937D7A0D0D33E47DCD6C84B312914B19C410A7A6D0E323177C5",
      INIT_02       =>
      X"C172B5A3D5B9C78DCDBBF5133194810CE3F4781CDD4ABDC529C497EFEB5553F8",
      INIT_03       =>
      X"0F68392934CC929E3769C51E095D22DEF25FA6BE20E3B20CCB7876DAD76E567C",
      INIT_04       =>
      X"07DFC62AEF1429601D3DEA5915AE4E65E3E079F9320922CD1C2D1F29C6F41430",
      INIT_05       =>
      X"06BBEA6BF06AD3C22D15E089DB669673E600343D102AF752C3C5C5A0E7B85767",
      INIT_06       =>
      X"32DFDD1509E1AF26C06A2A131B718699086EF9842AB062860DB5918616DA7878",
      INIT_07       =>
      X"E9233A7FE4A7FCF3DA0C1670E22F2650153FC3CAE53F83D3EAC56132CBE2A0EC",
      INIT_08       =>
      X"DBA7617FD3C74A273C17DDD833EF0A190BE783FE0D03B478D6B11FC036393599",
      INIT_09       =>
      X"E7E29A79220024553212697D11082202DB4439EB01A795BC23F241793FDDA378",
      INIT_0A       =>
      X"18FD51DACE195EB1FA3343230D1AB0EEDB39819C305193FD0CB086DBFFC7FB03",
      INIT_0B       =>
      X"039E2E8DF04B052312E512960D64F8F4C727CAA4EE3D15A4F358E28424F8A455",
      INIT_0C       =>
      X"39443AEA392C9DEDE34CFCB1396697731D853C6ECF85B28A3D4EB99B29963256",
      INIT_0D       =>
      X"2CAE9829C029FAA53688992AECE69D261847602CD48874D5FAD433A9C73F3E2A",
      INIT_0E       =>
      X"CFA77618295122CCD6017876EAAED1C4D053D0F2C7E819C5307B8EA103392005",
      INIT_0F       =>
      X"14097D5B1A5D8279071A45DF2A734B05D6BF53EDD6CF40BCD78E386F095A5AF9" )
    port map (ADDR  => addrE,
              CLK   => clk,
              DI    => x"00000000",
              DIP   => x"0",
              EN    => '1',
              SSR   => '0',
              WE    => '0',
              DO    => doE,
              DOP   => open);

  MEM_F : RAMB16_S36
    generic map (
      INIT_00       =>
      X"D46F6FDEF713D1D7EABB57B6CD3031B4FDCF96EDF18EB9C929E335030468FF7A",
      INIT_01       =>
      X"C55DFFD93F24C0AC2CE0CAAE0224DFD5D27628842CB6D00A0B9C46AB258F8B5E",
      INIT_02       =>
      X"2668ADDFD7B2A12B3F02F397DD0E52E6C80B2B13D5B1D0CBC70CDA711D5C594F",
      INIT_03       =>
      X"FA052740150DF46517858445359C27C6C104770B3D2801CCEE81E1E7D6912C06",
      INIT_04       =>
      X"D6E7914123085ADAEEE89003F15805E30E98EAFC37D4BE2CC69CAE2E0168B948",
      INIT_05       =>
      X"D9FC4EE00207B65BE8827A71FC9FF591FCA9B682E95DB9C50FBF2AE33A84D6AE",
      INIT_06       =>
      X"2D4DA6C2F30655A6F9BA1B1D16BC7ABD0C9DA7C7E20779F317B98726EF8F54E1",
      INIT_07       =>
      X"091C94FED7DD4C0903601232C7B3DBB61DD824C92E521DCDF02E5772283BFD04",
      INIT_08       =>
      X"F91F70E5D23C57833ABDDAD3FE9A9A373B54C642D7B57FF9CFB20A3509FCC05F",
      INIT_09       =>
      X"D3ABE099E1194A27F7D0DDC2241C8BB8C71CFB4735C92767FB9A11480A7D05B6",
      INIT_0A       =>
      X"2516DC3A13948666D34FDE063CDADF362646DFA4204988600320C419CF8A64E8",
      INIT_0B       =>
      X"0F4376C3D44EA62B1ACC4D0BC546B6640B32112E02EF010301E6A433037E3578",
      INIT_0C       =>
      X"313F06AC2238625B1CD49488E6C200F7E918F1770A983D05EC0426242A7E5740",
      INIT_0D       =>
      X"DF5CCC6BD0371221D9754C19CFD267833C8B3188385C01F3180189C2D86EA5D0",
      INIT_0E       =>
      X"074EADFEFE87CBA219383275C3D078871970EF68C5A3AC0F30809A811C961032",
      INIT_0F       =>
      X"06C170EF2FA903CEE6CF65571C4319AFE0658D0BD280BF2CC176CCA4DB1ED6A7" )
    port map (ADDR  => addrF,
              CLK   => clk,
              DI    => x"00000000",
              DIP   => x"0",
              EN    => '1',
              SSR   => '0',
              WE    => '0',
              DO    => doF,
              DOP   => open);

end GENERATED;
